module ALU_Reg (A_Mux_input, B_Mux_input, clk, decoder_input);
input [3:0] A_Mux_input, B_Mux_input, decoder_input; 


endmodule 